

module PC_Adder (a,b,c);

    input [31:0]a,b;
    output [31:0]c;

    assign c = a + b;
    
endmodule // add the 32 bit mer=iry address of one point to another point to get to specifed location for PC